/****************************************************************************
 * execution_stage.sv
 ****************************************************************************/
`include "integer.sv"

/**
 * Module: Execution_Stage
 * 
 * TODO: Add module documentation
 */
module Execution_Stage(input next);

Integer_Unit integer_unit(next);

/* TODO: Floating Point Unit */

endmodule
