`include "defines.sv"


module L1_DCache();
	
	
endmodule