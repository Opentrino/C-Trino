/****************************************************************************
 * l3_cache.sv
 ****************************************************************************/

/**
 * Module: L3_Cache
 * 
 * TODO: Add module documentation
 */
module L3_Cache(input next);


endmodule


