/****************************************************************************
 * memory_access_stage.sv
 ****************************************************************************/

/**
 * Module: Memory_Access_Stage
 * 
 * TODO: Add module documentation
 */
module Memory_Access_Stage(input next);

/* TODO: Implement Load and Store */
	
endmodule
