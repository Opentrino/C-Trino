/****************************************************************************
 * register_file.sv
 ****************************************************************************/

/**
 * Module: RegFile
 * 
 * TODO: Add module documentation
 */
module RegFile(input next);


endmodule
