`include "defines.sv"

module L2_Cache(input next);
	always@(next) begin 
		
	end
endmodule