`include "defines.sv"


module L1_DCache(input next);
	always@(next) begin
		
	end
endmodule