/****************************************************************************
 * predecode_stage.sv
 ****************************************************************************/

/**
 * Module: Stage_PreDecode
 * 
 * TODO: Add module documentation
 */
module Stage_PreDecode(input next);


endmodule
