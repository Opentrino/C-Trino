`ifndef DEFINES_SV_
`define DEFINES_SV_

/**********************/
/* MEMORY RAM DEFINES */
/**********************/
`define MEMORY_SIZE 256
`define MEMORY_WIDTH 8
`define MEMORY_SIZE_ENC ($clog2(`MEMORY_SIZE) - 1)
/**********************/

/*****************************/
/* 1: PREFETCH STAGE DEFINES */
/*****************************/

/*****************************/
	
/******************************/
/* 2: PREDECODE STAGE DEFINES */
/******************************/

/******************************/
	
/******************************/
/* 3: MICROCODE STAGE DEFINES */
/******************************/
`define UC_CTRL_WIDTH 32
`define UC_FUNC_WIDTH 32
`define UC_CTRL_DEPTH 200
`define UC_SEGMENT_MAXCOUNT 200
`define UC_CALLSTACK_SIZE 256
/******************************/

/***********************************/
/* 4: RENAME/REORDER STAGE DEFINES */
/***********************************/

/***********************************/

/**************************/
/* 5: ISSUE STAGE DEFINES */
/**************************/

/**************************/

/****************************/
/* 6: EXECUTE STAGE DEFINES */
/****************************/

/****************************/
	
/**********************************/
/* 7: MEMORY ACCESS STAGE DEFINES */
/**********************************/

/**********************************/

/******************************/
/* 8: WRITEBACK STAGE DEFINES */
/******************************/

/******************************/

/***************************/
/* 9: COMMIT STAGE DEFINES */
/***************************/

/***************************/

/********************************/
/* L1 INSTRUCTION CACHE DEFINES */
/********************************/

/********************************/

/*************************/
/* L1 DATA CACHE DEFINES */
/*************************/

/*************************/	

/********************/
/* L2 CACHE DEFINES */
/********************/

/********************/

/********************/
/* L3 CACHE DEFINES */
/********************/

/********************/

/******************/
/* UNCORE DEFINES */
/******************/

/******************/

`endif