module  name(rst,clk);
input rst;
input clk;

endmodule
