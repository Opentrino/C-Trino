`include "defines.sv"

module L2_Cache();
	
	
endmodule