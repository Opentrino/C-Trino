`include "defines.sv"


module L1_ICache();
	
	
endmodule