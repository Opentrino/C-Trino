`include "defines.sv"

/*
 ********************************************
 * 1- Fetch Stage
 *  1.1- Next Fetch Address prediction
 *    1.1.1- Branch Target Buffer (BTB)
 *    1.1.2- Next Sequential Fetch addr
 *    1.1.3- Branch Predictor
 *    1.1.4- Return Address Stack (RAS)
 *  1.2- Fetch address calculation
 *    1.2.1- Calculate address tag + index + offset
 *  1.3- ICache Access
 *    1.3.1- ICache Data Array
 *    1.3.2- ICache Tag Array
 *    1.3.3- ITLB Array
 *  1.4- Instruction drive to decode stage
 *    1.4.1- Aligner
 ********************************************
 */

/* STEPS: 
 * 
 */

module Stage_Fetch();
	

endmodule