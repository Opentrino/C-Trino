`include "defines.sv"

module L1_ICache(input next);
	always@(next) begin
		
	end
endmodule