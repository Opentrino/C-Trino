module core_main;

endmodule